`timescale 1ns/1ns
`include "axi4_lite.svh"

module topTB();

endmodule