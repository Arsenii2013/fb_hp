//`define PCIE_PIPE_STACK